magic
tech gf180mcuD
magscale 1 5
timestamp 1701413170
<< obsm1 >>
rect 672 855 149296 148206
<< metal2 >>
rect 7728 0 7784 400
rect 8176 0 8232 400
rect 8624 0 8680 400
rect 9072 0 9128 400
rect 9520 0 9576 400
rect 9968 0 10024 400
rect 10416 0 10472 400
rect 10864 0 10920 400
rect 11312 0 11368 400
rect 11760 0 11816 400
rect 12208 0 12264 400
rect 12656 0 12712 400
rect 13104 0 13160 400
rect 13552 0 13608 400
rect 14000 0 14056 400
rect 14448 0 14504 400
rect 14896 0 14952 400
rect 15344 0 15400 400
rect 15792 0 15848 400
rect 16240 0 16296 400
rect 16688 0 16744 400
rect 17136 0 17192 400
rect 17584 0 17640 400
rect 18032 0 18088 400
rect 18480 0 18536 400
rect 18928 0 18984 400
rect 19376 0 19432 400
rect 19824 0 19880 400
rect 20272 0 20328 400
rect 20720 0 20776 400
rect 21168 0 21224 400
rect 21616 0 21672 400
rect 22064 0 22120 400
rect 22512 0 22568 400
rect 22960 0 23016 400
rect 23408 0 23464 400
rect 23856 0 23912 400
rect 24304 0 24360 400
rect 24752 0 24808 400
rect 25200 0 25256 400
rect 25648 0 25704 400
rect 26096 0 26152 400
rect 26544 0 26600 400
rect 26992 0 27048 400
rect 27440 0 27496 400
rect 27888 0 27944 400
rect 28336 0 28392 400
rect 28784 0 28840 400
rect 29232 0 29288 400
rect 29680 0 29736 400
rect 30128 0 30184 400
rect 30576 0 30632 400
rect 31024 0 31080 400
rect 31472 0 31528 400
rect 31920 0 31976 400
rect 32368 0 32424 400
rect 32816 0 32872 400
rect 33264 0 33320 400
rect 33712 0 33768 400
rect 34160 0 34216 400
rect 34608 0 34664 400
rect 35056 0 35112 400
rect 35504 0 35560 400
rect 35952 0 36008 400
rect 36400 0 36456 400
rect 36848 0 36904 400
rect 37296 0 37352 400
rect 37744 0 37800 400
rect 38192 0 38248 400
rect 38640 0 38696 400
rect 39088 0 39144 400
rect 39536 0 39592 400
rect 39984 0 40040 400
rect 40432 0 40488 400
rect 40880 0 40936 400
rect 41328 0 41384 400
rect 41776 0 41832 400
rect 42224 0 42280 400
rect 42672 0 42728 400
rect 43120 0 43176 400
rect 43568 0 43624 400
rect 44016 0 44072 400
rect 44464 0 44520 400
rect 44912 0 44968 400
rect 45360 0 45416 400
rect 45808 0 45864 400
rect 46256 0 46312 400
rect 46704 0 46760 400
rect 47152 0 47208 400
rect 47600 0 47656 400
rect 48048 0 48104 400
rect 48496 0 48552 400
rect 48944 0 49000 400
rect 49392 0 49448 400
rect 49840 0 49896 400
rect 50288 0 50344 400
rect 50736 0 50792 400
rect 51184 0 51240 400
rect 51632 0 51688 400
rect 52080 0 52136 400
rect 52528 0 52584 400
rect 52976 0 53032 400
rect 53424 0 53480 400
rect 53872 0 53928 400
rect 54320 0 54376 400
rect 54768 0 54824 400
rect 55216 0 55272 400
rect 55664 0 55720 400
rect 56112 0 56168 400
rect 56560 0 56616 400
rect 57008 0 57064 400
rect 57456 0 57512 400
rect 57904 0 57960 400
rect 58352 0 58408 400
rect 58800 0 58856 400
rect 59248 0 59304 400
rect 59696 0 59752 400
rect 60144 0 60200 400
rect 60592 0 60648 400
rect 61040 0 61096 400
rect 61488 0 61544 400
rect 61936 0 61992 400
rect 62384 0 62440 400
rect 62832 0 62888 400
rect 63280 0 63336 400
rect 63728 0 63784 400
rect 64176 0 64232 400
rect 64624 0 64680 400
rect 65072 0 65128 400
rect 65520 0 65576 400
rect 65968 0 66024 400
rect 66416 0 66472 400
rect 66864 0 66920 400
rect 67312 0 67368 400
rect 67760 0 67816 400
rect 68208 0 68264 400
rect 68656 0 68712 400
rect 69104 0 69160 400
rect 69552 0 69608 400
rect 70000 0 70056 400
rect 70448 0 70504 400
rect 70896 0 70952 400
rect 71344 0 71400 400
rect 71792 0 71848 400
rect 72240 0 72296 400
rect 72688 0 72744 400
rect 73136 0 73192 400
rect 73584 0 73640 400
rect 74032 0 74088 400
rect 74480 0 74536 400
rect 74928 0 74984 400
rect 75376 0 75432 400
rect 75824 0 75880 400
rect 76272 0 76328 400
rect 76720 0 76776 400
rect 77168 0 77224 400
rect 77616 0 77672 400
rect 78064 0 78120 400
rect 78512 0 78568 400
rect 78960 0 79016 400
rect 79408 0 79464 400
rect 79856 0 79912 400
rect 80304 0 80360 400
rect 80752 0 80808 400
rect 81200 0 81256 400
rect 81648 0 81704 400
rect 82096 0 82152 400
rect 82544 0 82600 400
rect 82992 0 83048 400
rect 83440 0 83496 400
rect 83888 0 83944 400
rect 84336 0 84392 400
rect 84784 0 84840 400
rect 85232 0 85288 400
rect 85680 0 85736 400
rect 86128 0 86184 400
rect 86576 0 86632 400
rect 87024 0 87080 400
rect 87472 0 87528 400
rect 87920 0 87976 400
rect 88368 0 88424 400
rect 88816 0 88872 400
rect 89264 0 89320 400
rect 89712 0 89768 400
rect 90160 0 90216 400
rect 90608 0 90664 400
rect 91056 0 91112 400
rect 91504 0 91560 400
rect 91952 0 92008 400
rect 92400 0 92456 400
rect 92848 0 92904 400
rect 93296 0 93352 400
rect 93744 0 93800 400
rect 94192 0 94248 400
rect 94640 0 94696 400
rect 95088 0 95144 400
rect 95536 0 95592 400
rect 95984 0 96040 400
rect 96432 0 96488 400
rect 96880 0 96936 400
rect 97328 0 97384 400
rect 97776 0 97832 400
rect 98224 0 98280 400
rect 98672 0 98728 400
rect 99120 0 99176 400
rect 99568 0 99624 400
rect 100016 0 100072 400
rect 100464 0 100520 400
rect 100912 0 100968 400
rect 101360 0 101416 400
rect 101808 0 101864 400
rect 102256 0 102312 400
rect 102704 0 102760 400
rect 103152 0 103208 400
rect 103600 0 103656 400
rect 104048 0 104104 400
rect 104496 0 104552 400
rect 104944 0 105000 400
rect 105392 0 105448 400
rect 105840 0 105896 400
rect 106288 0 106344 400
rect 106736 0 106792 400
rect 107184 0 107240 400
rect 107632 0 107688 400
rect 108080 0 108136 400
rect 108528 0 108584 400
rect 108976 0 109032 400
rect 109424 0 109480 400
rect 109872 0 109928 400
rect 110320 0 110376 400
rect 110768 0 110824 400
rect 111216 0 111272 400
rect 111664 0 111720 400
rect 112112 0 112168 400
rect 112560 0 112616 400
rect 113008 0 113064 400
rect 113456 0 113512 400
rect 113904 0 113960 400
rect 114352 0 114408 400
rect 114800 0 114856 400
rect 115248 0 115304 400
rect 115696 0 115752 400
rect 116144 0 116200 400
rect 116592 0 116648 400
rect 117040 0 117096 400
rect 117488 0 117544 400
rect 117936 0 117992 400
rect 118384 0 118440 400
rect 118832 0 118888 400
rect 119280 0 119336 400
rect 119728 0 119784 400
rect 120176 0 120232 400
rect 120624 0 120680 400
rect 121072 0 121128 400
rect 121520 0 121576 400
rect 121968 0 122024 400
rect 122416 0 122472 400
rect 122864 0 122920 400
rect 123312 0 123368 400
rect 123760 0 123816 400
rect 124208 0 124264 400
rect 124656 0 124712 400
rect 125104 0 125160 400
rect 125552 0 125608 400
rect 126000 0 126056 400
rect 126448 0 126504 400
rect 126896 0 126952 400
rect 127344 0 127400 400
rect 127792 0 127848 400
rect 128240 0 128296 400
rect 128688 0 128744 400
rect 129136 0 129192 400
rect 129584 0 129640 400
rect 130032 0 130088 400
rect 130480 0 130536 400
rect 130928 0 130984 400
rect 131376 0 131432 400
rect 131824 0 131880 400
rect 132272 0 132328 400
rect 132720 0 132776 400
rect 133168 0 133224 400
rect 133616 0 133672 400
rect 134064 0 134120 400
rect 134512 0 134568 400
rect 134960 0 135016 400
rect 135408 0 135464 400
rect 135856 0 135912 400
rect 136304 0 136360 400
rect 136752 0 136808 400
rect 137200 0 137256 400
rect 137648 0 137704 400
rect 138096 0 138152 400
rect 138544 0 138600 400
rect 138992 0 139048 400
rect 139440 0 139496 400
rect 139888 0 139944 400
rect 140336 0 140392 400
rect 140784 0 140840 400
rect 141232 0 141288 400
rect 141680 0 141736 400
rect 142128 0 142184 400
<< obsm2 >>
rect 854 430 149114 148195
rect 854 350 7698 430
rect 7814 350 8146 430
rect 8262 350 8594 430
rect 8710 350 9042 430
rect 9158 350 9490 430
rect 9606 350 9938 430
rect 10054 350 10386 430
rect 10502 350 10834 430
rect 10950 350 11282 430
rect 11398 350 11730 430
rect 11846 350 12178 430
rect 12294 350 12626 430
rect 12742 350 13074 430
rect 13190 350 13522 430
rect 13638 350 13970 430
rect 14086 350 14418 430
rect 14534 350 14866 430
rect 14982 350 15314 430
rect 15430 350 15762 430
rect 15878 350 16210 430
rect 16326 350 16658 430
rect 16774 350 17106 430
rect 17222 350 17554 430
rect 17670 350 18002 430
rect 18118 350 18450 430
rect 18566 350 18898 430
rect 19014 350 19346 430
rect 19462 350 19794 430
rect 19910 350 20242 430
rect 20358 350 20690 430
rect 20806 350 21138 430
rect 21254 350 21586 430
rect 21702 350 22034 430
rect 22150 350 22482 430
rect 22598 350 22930 430
rect 23046 350 23378 430
rect 23494 350 23826 430
rect 23942 350 24274 430
rect 24390 350 24722 430
rect 24838 350 25170 430
rect 25286 350 25618 430
rect 25734 350 26066 430
rect 26182 350 26514 430
rect 26630 350 26962 430
rect 27078 350 27410 430
rect 27526 350 27858 430
rect 27974 350 28306 430
rect 28422 350 28754 430
rect 28870 350 29202 430
rect 29318 350 29650 430
rect 29766 350 30098 430
rect 30214 350 30546 430
rect 30662 350 30994 430
rect 31110 350 31442 430
rect 31558 350 31890 430
rect 32006 350 32338 430
rect 32454 350 32786 430
rect 32902 350 33234 430
rect 33350 350 33682 430
rect 33798 350 34130 430
rect 34246 350 34578 430
rect 34694 350 35026 430
rect 35142 350 35474 430
rect 35590 350 35922 430
rect 36038 350 36370 430
rect 36486 350 36818 430
rect 36934 350 37266 430
rect 37382 350 37714 430
rect 37830 350 38162 430
rect 38278 350 38610 430
rect 38726 350 39058 430
rect 39174 350 39506 430
rect 39622 350 39954 430
rect 40070 350 40402 430
rect 40518 350 40850 430
rect 40966 350 41298 430
rect 41414 350 41746 430
rect 41862 350 42194 430
rect 42310 350 42642 430
rect 42758 350 43090 430
rect 43206 350 43538 430
rect 43654 350 43986 430
rect 44102 350 44434 430
rect 44550 350 44882 430
rect 44998 350 45330 430
rect 45446 350 45778 430
rect 45894 350 46226 430
rect 46342 350 46674 430
rect 46790 350 47122 430
rect 47238 350 47570 430
rect 47686 350 48018 430
rect 48134 350 48466 430
rect 48582 350 48914 430
rect 49030 350 49362 430
rect 49478 350 49810 430
rect 49926 350 50258 430
rect 50374 350 50706 430
rect 50822 350 51154 430
rect 51270 350 51602 430
rect 51718 350 52050 430
rect 52166 350 52498 430
rect 52614 350 52946 430
rect 53062 350 53394 430
rect 53510 350 53842 430
rect 53958 350 54290 430
rect 54406 350 54738 430
rect 54854 350 55186 430
rect 55302 350 55634 430
rect 55750 350 56082 430
rect 56198 350 56530 430
rect 56646 350 56978 430
rect 57094 350 57426 430
rect 57542 350 57874 430
rect 57990 350 58322 430
rect 58438 350 58770 430
rect 58886 350 59218 430
rect 59334 350 59666 430
rect 59782 350 60114 430
rect 60230 350 60562 430
rect 60678 350 61010 430
rect 61126 350 61458 430
rect 61574 350 61906 430
rect 62022 350 62354 430
rect 62470 350 62802 430
rect 62918 350 63250 430
rect 63366 350 63698 430
rect 63814 350 64146 430
rect 64262 350 64594 430
rect 64710 350 65042 430
rect 65158 350 65490 430
rect 65606 350 65938 430
rect 66054 350 66386 430
rect 66502 350 66834 430
rect 66950 350 67282 430
rect 67398 350 67730 430
rect 67846 350 68178 430
rect 68294 350 68626 430
rect 68742 350 69074 430
rect 69190 350 69522 430
rect 69638 350 69970 430
rect 70086 350 70418 430
rect 70534 350 70866 430
rect 70982 350 71314 430
rect 71430 350 71762 430
rect 71878 350 72210 430
rect 72326 350 72658 430
rect 72774 350 73106 430
rect 73222 350 73554 430
rect 73670 350 74002 430
rect 74118 350 74450 430
rect 74566 350 74898 430
rect 75014 350 75346 430
rect 75462 350 75794 430
rect 75910 350 76242 430
rect 76358 350 76690 430
rect 76806 350 77138 430
rect 77254 350 77586 430
rect 77702 350 78034 430
rect 78150 350 78482 430
rect 78598 350 78930 430
rect 79046 350 79378 430
rect 79494 350 79826 430
rect 79942 350 80274 430
rect 80390 350 80722 430
rect 80838 350 81170 430
rect 81286 350 81618 430
rect 81734 350 82066 430
rect 82182 350 82514 430
rect 82630 350 82962 430
rect 83078 350 83410 430
rect 83526 350 83858 430
rect 83974 350 84306 430
rect 84422 350 84754 430
rect 84870 350 85202 430
rect 85318 350 85650 430
rect 85766 350 86098 430
rect 86214 350 86546 430
rect 86662 350 86994 430
rect 87110 350 87442 430
rect 87558 350 87890 430
rect 88006 350 88338 430
rect 88454 350 88786 430
rect 88902 350 89234 430
rect 89350 350 89682 430
rect 89798 350 90130 430
rect 90246 350 90578 430
rect 90694 350 91026 430
rect 91142 350 91474 430
rect 91590 350 91922 430
rect 92038 350 92370 430
rect 92486 350 92818 430
rect 92934 350 93266 430
rect 93382 350 93714 430
rect 93830 350 94162 430
rect 94278 350 94610 430
rect 94726 350 95058 430
rect 95174 350 95506 430
rect 95622 350 95954 430
rect 96070 350 96402 430
rect 96518 350 96850 430
rect 96966 350 97298 430
rect 97414 350 97746 430
rect 97862 350 98194 430
rect 98310 350 98642 430
rect 98758 350 99090 430
rect 99206 350 99538 430
rect 99654 350 99986 430
rect 100102 350 100434 430
rect 100550 350 100882 430
rect 100998 350 101330 430
rect 101446 350 101778 430
rect 101894 350 102226 430
rect 102342 350 102674 430
rect 102790 350 103122 430
rect 103238 350 103570 430
rect 103686 350 104018 430
rect 104134 350 104466 430
rect 104582 350 104914 430
rect 105030 350 105362 430
rect 105478 350 105810 430
rect 105926 350 106258 430
rect 106374 350 106706 430
rect 106822 350 107154 430
rect 107270 350 107602 430
rect 107718 350 108050 430
rect 108166 350 108498 430
rect 108614 350 108946 430
rect 109062 350 109394 430
rect 109510 350 109842 430
rect 109958 350 110290 430
rect 110406 350 110738 430
rect 110854 350 111186 430
rect 111302 350 111634 430
rect 111750 350 112082 430
rect 112198 350 112530 430
rect 112646 350 112978 430
rect 113094 350 113426 430
rect 113542 350 113874 430
rect 113990 350 114322 430
rect 114438 350 114770 430
rect 114886 350 115218 430
rect 115334 350 115666 430
rect 115782 350 116114 430
rect 116230 350 116562 430
rect 116678 350 117010 430
rect 117126 350 117458 430
rect 117574 350 117906 430
rect 118022 350 118354 430
rect 118470 350 118802 430
rect 118918 350 119250 430
rect 119366 350 119698 430
rect 119814 350 120146 430
rect 120262 350 120594 430
rect 120710 350 121042 430
rect 121158 350 121490 430
rect 121606 350 121938 430
rect 122054 350 122386 430
rect 122502 350 122834 430
rect 122950 350 123282 430
rect 123398 350 123730 430
rect 123846 350 124178 430
rect 124294 350 124626 430
rect 124742 350 125074 430
rect 125190 350 125522 430
rect 125638 350 125970 430
rect 126086 350 126418 430
rect 126534 350 126866 430
rect 126982 350 127314 430
rect 127430 350 127762 430
rect 127878 350 128210 430
rect 128326 350 128658 430
rect 128774 350 129106 430
rect 129222 350 129554 430
rect 129670 350 130002 430
rect 130118 350 130450 430
rect 130566 350 130898 430
rect 131014 350 131346 430
rect 131462 350 131794 430
rect 131910 350 132242 430
rect 132358 350 132690 430
rect 132806 350 133138 430
rect 133254 350 133586 430
rect 133702 350 134034 430
rect 134150 350 134482 430
rect 134598 350 134930 430
rect 135046 350 135378 430
rect 135494 350 135826 430
rect 135942 350 136274 430
rect 136390 350 136722 430
rect 136838 350 137170 430
rect 137286 350 137618 430
rect 137734 350 138066 430
rect 138182 350 138514 430
rect 138630 350 138962 430
rect 139078 350 139410 430
rect 139526 350 139858 430
rect 139974 350 140306 430
rect 140422 350 140754 430
rect 140870 350 141202 430
rect 141318 350 141650 430
rect 141766 350 142098 430
rect 142214 350 149114 430
<< metal3 >>
rect 0 145712 400 145768
rect 149600 145712 150000 145768
rect 0 139552 400 139608
rect 149600 139552 150000 139608
rect 0 133392 400 133448
rect 149600 133392 150000 133448
rect 0 127232 400 127288
rect 149600 127232 150000 127288
rect 0 121072 400 121128
rect 149600 121072 150000 121128
rect 0 114912 400 114968
rect 149600 114912 150000 114968
rect 0 108752 400 108808
rect 149600 108752 150000 108808
rect 0 102592 400 102648
rect 149600 102592 150000 102648
rect 0 96432 400 96488
rect 149600 96432 150000 96488
rect 0 90272 400 90328
rect 149600 90272 150000 90328
rect 0 84112 400 84168
rect 149600 84112 150000 84168
rect 0 77952 400 78008
rect 149600 77952 150000 78008
rect 0 71792 400 71848
rect 149600 71792 150000 71848
rect 0 65632 400 65688
rect 149600 65632 150000 65688
rect 0 59472 400 59528
rect 149600 59472 150000 59528
rect 0 53312 400 53368
rect 149600 53312 150000 53368
rect 0 47152 400 47208
rect 149600 47152 150000 47208
rect 0 40992 400 41048
rect 149600 40992 150000 41048
rect 0 34832 400 34888
rect 149600 34832 150000 34888
rect 0 28672 400 28728
rect 149600 28672 150000 28728
rect 0 22512 400 22568
rect 149600 22512 150000 22568
rect 0 16352 400 16408
rect 149600 16352 150000 16408
rect 0 10192 400 10248
rect 149600 10192 150000 10248
rect 0 4032 400 4088
rect 149600 4032 150000 4088
<< obsm3 >>
rect 400 145798 149600 148190
rect 430 145682 149570 145798
rect 400 139638 149600 145682
rect 430 139522 149570 139638
rect 400 133478 149600 139522
rect 430 133362 149570 133478
rect 400 127318 149600 133362
rect 430 127202 149570 127318
rect 400 121158 149600 127202
rect 430 121042 149570 121158
rect 400 114998 149600 121042
rect 430 114882 149570 114998
rect 400 108838 149600 114882
rect 430 108722 149570 108838
rect 400 102678 149600 108722
rect 430 102562 149570 102678
rect 400 96518 149600 102562
rect 430 96402 149570 96518
rect 400 90358 149600 96402
rect 430 90242 149570 90358
rect 400 84198 149600 90242
rect 430 84082 149570 84198
rect 400 78038 149600 84082
rect 430 77922 149570 78038
rect 400 71878 149600 77922
rect 430 71762 149570 71878
rect 400 65718 149600 71762
rect 430 65602 149570 65718
rect 400 59558 149600 65602
rect 430 59442 149570 59558
rect 400 53398 149600 59442
rect 430 53282 149570 53398
rect 400 47238 149600 53282
rect 430 47122 149570 47238
rect 400 41078 149600 47122
rect 430 40962 149570 41078
rect 400 34918 149600 40962
rect 430 34802 149570 34918
rect 400 28758 149600 34802
rect 430 28642 149570 28758
rect 400 22598 149600 28642
rect 430 22482 149570 22598
rect 400 16438 149600 22482
rect 430 16322 149570 16438
rect 400 10278 149600 16322
rect 430 10162 149570 10278
rect 400 4118 149600 10162
rect 430 4002 149570 4118
rect 400 1554 149600 4002
<< metal4 >>
rect 2224 1538 2384 148206
rect 9904 1538 10064 148206
rect 17584 1538 17744 148206
rect 25264 1538 25424 148206
rect 32944 1538 33104 148206
rect 40624 1538 40784 148206
rect 48304 1538 48464 148206
rect 55984 1538 56144 148206
rect 63664 1538 63824 148206
rect 71344 1538 71504 148206
rect 79024 1538 79184 148206
rect 86704 1538 86864 148206
rect 94384 1538 94544 148206
rect 102064 1538 102224 148206
rect 109744 1538 109904 148206
rect 117424 1538 117584 148206
rect 125104 1538 125264 148206
rect 132784 1538 132944 148206
rect 140464 1538 140624 148206
rect 148144 1538 148304 148206
<< obsm4 >>
rect 5838 3313 9874 120335
rect 10094 3313 17554 120335
rect 17774 3313 25234 120335
rect 25454 3313 32914 120335
rect 33134 3313 40594 120335
rect 40814 3313 48274 120335
rect 48494 3313 55954 120335
rect 56174 3313 63634 120335
rect 63854 3313 71314 120335
rect 71534 3313 78994 120335
rect 79214 3313 86674 120335
rect 86894 3313 94354 120335
rect 94574 3313 102034 120335
rect 102254 3313 109714 120335
rect 109934 3313 117394 120335
rect 117614 3313 125074 120335
rect 125294 3313 132754 120335
rect 132974 3313 140434 120335
rect 140654 3313 142338 120335
<< labels >>
rlabel metal3 s 149600 4032 150000 4088 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 108752 400 108808 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 90272 400 90328 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 71792 400 71848 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 53312 400 53368 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 34832 400 34888 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 16352 400 16408 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 149600 22512 150000 22568 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 149600 40992 150000 41048 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 149600 59472 150000 59528 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 149600 77952 150000 78008 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 149600 96432 150000 96488 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 149600 114912 150000 114968 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 149600 133392 150000 133448 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 145712 400 145768 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 127232 400 127288 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 149600 16352 150000 16408 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 96432 400 96488 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 77952 400 78008 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 59472 400 59528 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 40992 400 41048 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 22512 400 22568 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 4032 400 4088 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 149600 34832 150000 34888 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 149600 53312 150000 53368 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 149600 71792 150000 71848 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 149600 90272 150000 90328 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 149600 108752 150000 108808 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 149600 127232 150000 127288 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 149600 145712 150000 145768 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 133392 400 133448 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 114912 400 114968 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 149600 10192 150000 10248 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 102592 400 102648 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 84112 400 84168 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 65632 400 65688 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 47152 400 47208 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 28672 400 28728 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 10192 400 10248 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 149600 28672 150000 28728 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 149600 47152 150000 47208 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 149600 65632 150000 65688 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 149600 84112 150000 84168 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 149600 102592 150000 102648 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 149600 121072 150000 121128 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 149600 139552 150000 139608 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 139552 400 139608 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 121072 400 121128 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 141232 0 141288 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 141680 0 141736 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 142128 0 142184 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 55216 0 55272 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 68656 0 68712 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 70000 0 70056 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 71344 0 71400 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 72688 0 72744 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 74032 0 74088 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 75376 0 75432 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 76720 0 76776 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 78064 0 78120 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 80752 0 80808 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 56560 0 56616 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 82096 0 82152 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 83440 0 83496 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 84784 0 84840 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 86128 0 86184 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 87472 0 87528 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 88816 0 88872 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 90160 0 90216 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 91504 0 91560 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 92848 0 92904 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 94192 0 94248 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 95536 0 95592 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 96880 0 96936 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 98224 0 98280 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 99568 0 99624 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 100912 0 100968 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 102256 0 102312 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 103600 0 103656 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 104944 0 105000 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 106288 0 106344 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 107632 0 107688 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 108976 0 109032 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 110320 0 110376 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 111664 0 111720 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 113008 0 113064 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 114352 0 114408 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 115696 0 115752 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 117040 0 117096 400 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 118384 0 118440 400 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 119728 0 119784 400 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 121072 0 121128 400 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 60592 0 60648 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 122416 0 122472 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 123760 0 123816 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 125104 0 125160 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 126448 0 126504 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 127792 0 127848 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 129136 0 129192 400 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 130480 0 130536 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 131824 0 131880 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 133168 0 133224 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 134512 0 134568 400 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 61936 0 61992 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 135856 0 135912 400 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 137200 0 137256 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 138544 0 138600 400 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 139888 0 139944 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 63280 0 63336 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 64624 0 64680 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 65968 0 66024 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 67312 0 67368 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 69104 0 69160 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 70448 0 70504 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 71792 0 71848 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 73136 0 73192 400 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 74480 0 74536 400 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 75824 0 75880 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 77168 0 77224 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 78512 0 78568 400 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 79856 0 79912 400 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 81200 0 81256 400 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 57008 0 57064 400 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 82544 0 82600 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 83888 0 83944 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 85232 0 85288 400 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 86576 0 86632 400 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 87920 0 87976 400 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 89264 0 89320 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 90608 0 90664 400 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 91952 0 92008 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 93296 0 93352 400 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 94640 0 94696 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 58352 0 58408 400 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 95984 0 96040 400 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 97328 0 97384 400 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 98672 0 98728 400 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 100016 0 100072 400 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 101360 0 101416 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 102704 0 102760 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 104048 0 104104 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 105392 0 105448 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 106736 0 106792 400 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 108080 0 108136 400 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 59696 0 59752 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 109424 0 109480 400 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 110768 0 110824 400 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 112112 0 112168 400 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 113456 0 113512 400 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 114800 0 114856 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 116144 0 116200 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 117488 0 117544 400 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 118832 0 118888 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 120176 0 120232 400 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 121520 0 121576 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 61040 0 61096 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 122864 0 122920 400 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 124208 0 124264 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 125552 0 125608 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 126896 0 126952 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 128240 0 128296 400 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 129584 0 129640 400 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 130928 0 130984 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 132272 0 132328 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 133616 0 133672 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 134960 0 135016 400 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 62384 0 62440 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 136304 0 136360 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 137648 0 137704 400 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 138992 0 139048 400 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 140336 0 140392 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 63728 0 63784 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 65072 0 65128 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 66416 0 66472 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 67760 0 67816 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 56112 0 56168 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 69552 0 69608 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 70896 0 70952 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 72240 0 72296 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 74928 0 74984 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 76272 0 76328 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 77616 0 77672 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 78960 0 79016 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 80304 0 80360 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 82992 0 83048 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 84336 0 84392 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 85680 0 85736 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 87024 0 87080 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 88368 0 88424 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 89712 0 89768 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 91056 0 91112 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 92400 0 92456 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 93744 0 93800 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 95088 0 95144 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 58800 0 58856 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 96432 0 96488 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 97776 0 97832 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 99120 0 99176 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 100464 0 100520 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 101808 0 101864 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 103152 0 103208 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 104496 0 104552 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 105840 0 105896 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 107184 0 107240 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 108528 0 108584 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 60144 0 60200 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 109872 0 109928 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 111216 0 111272 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 112560 0 112616 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 113904 0 113960 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 115248 0 115304 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 116592 0 116648 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 117936 0 117992 400 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 119280 0 119336 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 120624 0 120680 400 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 121968 0 122024 400 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 61488 0 61544 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 123312 0 123368 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 124656 0 124712 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 126000 0 126056 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 127344 0 127400 400 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 128688 0 128744 400 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 130032 0 130088 400 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 131376 0 131432 400 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 132720 0 132776 400 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 134064 0 134120 400 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 62832 0 62888 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 136752 0 136808 400 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 138096 0 138152 400 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 139440 0 139496 400 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 140784 0 140840 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 64176 0 64232 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 65520 0 65576 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 66864 0 66920 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal4 s 2224 1538 2384 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 148206 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 148206 6 vss
port 245 nsew ground bidirectional
rlabel metal2 s 7728 0 7784 400 6 wb_clk_i
port 246 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wb_rst_i
port 247 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 wbs_ack_o
port 248 nsew signal output
rlabel metal2 s 10416 0 10472 400 6 wbs_adr_i[0]
port 249 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 wbs_adr_i[10]
port 250 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 wbs_adr_i[11]
port 251 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 wbs_adr_i[12]
port 252 nsew signal input
rlabel metal2 s 29680 0 29736 400 6 wbs_adr_i[13]
port 253 nsew signal input
rlabel metal2 s 31024 0 31080 400 6 wbs_adr_i[14]
port 254 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 wbs_adr_i[15]
port 255 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 wbs_adr_i[16]
port 256 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 wbs_adr_i[17]
port 257 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 wbs_adr_i[18]
port 258 nsew signal input
rlabel metal2 s 37744 0 37800 400 6 wbs_adr_i[19]
port 259 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_adr_i[1]
port 260 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 wbs_adr_i[20]
port 261 nsew signal input
rlabel metal2 s 40432 0 40488 400 6 wbs_adr_i[21]
port 262 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 wbs_adr_i[22]
port 263 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 wbs_adr_i[23]
port 264 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 wbs_adr_i[24]
port 265 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 wbs_adr_i[25]
port 266 nsew signal input
rlabel metal2 s 47152 0 47208 400 6 wbs_adr_i[26]
port 267 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 wbs_adr_i[27]
port 268 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 wbs_adr_i[28]
port 269 nsew signal input
rlabel metal2 s 51184 0 51240 400 6 wbs_adr_i[29]
port 270 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 wbs_adr_i[2]
port 271 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 wbs_adr_i[30]
port 272 nsew signal input
rlabel metal2 s 53872 0 53928 400 6 wbs_adr_i[31]
port 273 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 wbs_adr_i[3]
port 274 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_adr_i[4]
port 275 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_adr_i[5]
port 276 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_adr_i[6]
port 277 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 wbs_adr_i[7]
port 278 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 wbs_adr_i[8]
port 279 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_adr_i[9]
port 280 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_cyc_i
port 281 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 wbs_dat_i[0]
port 282 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 wbs_dat_i[10]
port 283 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_dat_i[11]
port 284 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_dat_i[12]
port 285 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 wbs_dat_i[13]
port 286 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 wbs_dat_i[14]
port 287 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 wbs_dat_i[15]
port 288 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 wbs_dat_i[16]
port 289 nsew signal input
rlabel metal2 s 35504 0 35560 400 6 wbs_dat_i[17]
port 290 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 wbs_dat_i[18]
port 291 nsew signal input
rlabel metal2 s 38192 0 38248 400 6 wbs_dat_i[19]
port 292 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 wbs_dat_i[1]
port 293 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 wbs_dat_i[20]
port 294 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 wbs_dat_i[21]
port 295 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 wbs_dat_i[22]
port 296 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 wbs_dat_i[23]
port 297 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 wbs_dat_i[24]
port 298 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 wbs_dat_i[25]
port 299 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 wbs_dat_i[26]
port 300 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 wbs_dat_i[27]
port 301 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 wbs_dat_i[28]
port 302 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 wbs_dat_i[29]
port 303 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_dat_i[2]
port 304 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 wbs_dat_i[30]
port 305 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 wbs_dat_i[31]
port 306 nsew signal input
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_i[3]
port 307 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 wbs_dat_i[4]
port 308 nsew signal input
rlabel metal2 s 19376 0 19432 400 6 wbs_dat_i[5]
port 309 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_dat_i[6]
port 310 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 wbs_dat_i[7]
port 311 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 wbs_dat_i[8]
port 312 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 wbs_dat_i[9]
port 313 nsew signal input
rlabel metal2 s 11312 0 11368 400 6 wbs_dat_o[0]
port 314 nsew signal output
rlabel metal2 s 26544 0 26600 400 6 wbs_dat_o[10]
port 315 nsew signal output
rlabel metal2 s 27888 0 27944 400 6 wbs_dat_o[11]
port 316 nsew signal output
rlabel metal2 s 29232 0 29288 400 6 wbs_dat_o[12]
port 317 nsew signal output
rlabel metal2 s 30576 0 30632 400 6 wbs_dat_o[13]
port 318 nsew signal output
rlabel metal2 s 31920 0 31976 400 6 wbs_dat_o[14]
port 319 nsew signal output
rlabel metal2 s 33264 0 33320 400 6 wbs_dat_o[15]
port 320 nsew signal output
rlabel metal2 s 34608 0 34664 400 6 wbs_dat_o[16]
port 321 nsew signal output
rlabel metal2 s 35952 0 36008 400 6 wbs_dat_o[17]
port 322 nsew signal output
rlabel metal2 s 37296 0 37352 400 6 wbs_dat_o[18]
port 323 nsew signal output
rlabel metal2 s 38640 0 38696 400 6 wbs_dat_o[19]
port 324 nsew signal output
rlabel metal2 s 13104 0 13160 400 6 wbs_dat_o[1]
port 325 nsew signal output
rlabel metal2 s 39984 0 40040 400 6 wbs_dat_o[20]
port 326 nsew signal output
rlabel metal2 s 41328 0 41384 400 6 wbs_dat_o[21]
port 327 nsew signal output
rlabel metal2 s 42672 0 42728 400 6 wbs_dat_o[22]
port 328 nsew signal output
rlabel metal2 s 44016 0 44072 400 6 wbs_dat_o[23]
port 329 nsew signal output
rlabel metal2 s 45360 0 45416 400 6 wbs_dat_o[24]
port 330 nsew signal output
rlabel metal2 s 46704 0 46760 400 6 wbs_dat_o[25]
port 331 nsew signal output
rlabel metal2 s 48048 0 48104 400 6 wbs_dat_o[26]
port 332 nsew signal output
rlabel metal2 s 49392 0 49448 400 6 wbs_dat_o[27]
port 333 nsew signal output
rlabel metal2 s 50736 0 50792 400 6 wbs_dat_o[28]
port 334 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 wbs_dat_o[29]
port 335 nsew signal output
rlabel metal2 s 14896 0 14952 400 6 wbs_dat_o[2]
port 336 nsew signal output
rlabel metal2 s 53424 0 53480 400 6 wbs_dat_o[30]
port 337 nsew signal output
rlabel metal2 s 54768 0 54824 400 6 wbs_dat_o[31]
port 338 nsew signal output
rlabel metal2 s 16688 0 16744 400 6 wbs_dat_o[3]
port 339 nsew signal output
rlabel metal2 s 18480 0 18536 400 6 wbs_dat_o[4]
port 340 nsew signal output
rlabel metal2 s 19824 0 19880 400 6 wbs_dat_o[5]
port 341 nsew signal output
rlabel metal2 s 21168 0 21224 400 6 wbs_dat_o[6]
port 342 nsew signal output
rlabel metal2 s 22512 0 22568 400 6 wbs_dat_o[7]
port 343 nsew signal output
rlabel metal2 s 23856 0 23912 400 6 wbs_dat_o[8]
port 344 nsew signal output
rlabel metal2 s 25200 0 25256 400 6 wbs_dat_o[9]
port 345 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 wbs_sel_i[0]
port 346 nsew signal input
rlabel metal2 s 13552 0 13608 400 6 wbs_sel_i[1]
port 347 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 wbs_sel_i[2]
port 348 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 wbs_sel_i[3]
port 349 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 wbs_stb_i
port 350 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_we_i
port 351 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 150000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35824808
string GDS_FILE /home/shahid/Desktop/test123/caravel_user_project/openlane/user_proj_example/runs/23_12_01_11_34/results/signoff/user_proj_example.magic.gds
string GDS_START 499170
<< end >>

